package brt_usb_seq_pkg;

`include "brt_uvm_methodology.svh"

import brt_usb_pkg::*;
import brt_usb_env_pkg::*;

`include "brt_usb_host_util_callback.sv"
`include "brt_usb_dev_util_callback.sv"
`include "brt_usb_xfer_seq_extends.sv"
`include "brt_usb_packet_seq_extends.sv"
`include "brt_usb_virtual_seq_extends.sv"

endpackage : brt_usb_seq_pkg
