interface brt_usb_if();
    brt_usb_20_serial_if brt_usb_20_serial_if();
    brt_usb_20_utmi_if   brt_usb_20_utmi_if();
    brt_usb_ss_serial_if brt_usb_ss_serial_if();

endinterface
