`include "brt_usb_base_virtual_sequence.sv"

// testcases
`include "brt_usb_all_test_sequence.sv"
