class brt_usb_multi_xfer_interleaving_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_multi_xfer_interleaving_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_multi_xfer_interleaving_vseq");
    super.new(name);
    //err_inject_cb = new();
  endfunction

  virtual task body();
    super.body();
    init_callback();
    //uvm_callbacks#(usb_protocol)::add(p_sequencer.agt.prot,err_inject_cb);
    p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[0].max_burst_size = 3;
    p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[1].max_burst_size = 3;
    p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[2].max_burst_size = 4;
    p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[5].max_burst_size = 1;
    p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[6].max_burst_size = 2;
    p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size = 2;
    p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size = 2;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    brt_usb_base_control_xfer_sequence ctrl_seq;

    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        begin
            bulk_out_xfer();
            bulk_out_xfer();
            bulk_out_xfer();
            bulk_out_xfer();
        end
        //// 2nd
        begin
            bulk_in_xfer();
            bulk_in_xfer();
            bulk_in_xfer();
            bulk_in_xfer();
        end
        // Interrupt
        begin
            interrupt_out_xfer();
            interrupt_out_xfer();
            interrupt_out_xfer();
            interrupt_out_xfer();
        end
        //// 2nd
        begin
            interrupt_in_xfer();
            interrupt_in_xfer();
            interrupt_in_xfer();
            interrupt_in_xfer();
        end
        // Iso
        begin
            isochronous_out_xfer();
            isochronous_out_xfer();
            isochronous_out_xfer();
            isochronous_out_xfer();
        end
        //// 2nd
        begin
            isochronous_in_xfer();
            isochronous_in_xfer();
            isochronous_in_xfer();
            isochronous_in_xfer();
        end
        // CTRL
        begin
            ctrl_xfer (.set_dir(0), .set_payload_size());
            ctrl_xfer (.set_dir(1), .set_payload_size());
            ctrl_xfer (.set_dir(0), .set_payload_size());
            ctrl_xfer (.set_dir(1), .set_payload_size());
        end
    join
  endtask
endclass

// Reset handshake
class brt_usb_reset_handshake_resume_vseq extends brt_usb_base_virtual_sequence;

  `brt_object_utils_begin(brt_usb_reset_handshake_resume_vseq)
  `brt_object_utils_end

  function new(string name="brt_usb_reset_handshake_resume_vseq");
    super.new(name);
  endfunction

  virtual task body();
    brt_usb_base_control_xfer_sequence              ctrl_seq;
    brt_usb_link_service_reset_sequence             reset_seq;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;
    brt_usb_agent_wait_for_link_usb_20_state_virtual_sequence wait_state;

    // Start
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::DEVICE_ATTACHED);
    // Reset device
    `brt_do_on(reset_seq, p_sequencer.link_service_sequencer) 

    `brt_info("DD", $sformatf("Wait for link state to ENABLE state"), UVM_LOW)
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    `brt_info("DD", $sformatf("link is ENABLE state"), UVM_LOW)

    #50us; 
    // reset 2nd time
    `brt_info("DD", $sformatf("link start to reset"), UVM_LOW)
    `brt_do_on(reset_seq, p_sequencer.link_service_sequencer) 
    `brt_info("DD", $sformatf("link is reseting"), UVM_LOW)
    // Wait ENABLE
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    `brt_info("DD", $sformatf("link is ENABLE state"), UVM_LOW)

    // let device enter suspend
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::SUSPENDED);

    #50us;
    // Host resume
    `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    #20us;

    init_callback();
    bulk_in_xfer();
    bulk_out_xfer();
    #10us;
  endtask
endclass

class brt_usb_reset_handshake_resume_w25_vseq extends brt_usb_base_virtual_sequence;

  `brt_object_utils_begin(brt_usb_reset_handshake_resume_w25_vseq)
  `brt_object_utils_end

  function new(string name="brt_usb_reset_handshake_resume_w25_vseq");
    super.new(name);
  endfunction

  virtual task body();
    brt_usb_base_control_xfer_sequence              ctrl_seq;
    brt_usb_link_service_reset_sequence             reset_seq;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;
    brt_usb_agent_wait_for_link_usb_20_state_virtual_sequence wait_state;

    super.body();
    host_cfg.tdchbit = 2.5us;

    // Start
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::DEVICE_ATTACHED);
    // Reset device
    `brt_do_on(reset_seq, p_sequencer.link_service_sequencer) 

    `brt_info("DD", $sformatf("Wait for link state to ENABLE state"), UVM_LOW)
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    `brt_info("DD", $sformatf("link is ENABLE state"), UVM_LOW)

    #50us; 
    // reset 2nd time
    `brt_info("DD", $sformatf("link start to reset"), UVM_LOW)
    `brt_do_on(reset_seq, p_sequencer.link_service_sequencer) 
    `brt_info("DD", $sformatf("link is reseting"), UVM_LOW)
    // Wait ENABLE
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    `brt_info("DD", $sformatf("link is ENABLE state"), UVM_LOW)

    // let device enter suspend
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::SUSPENDED);

    #50us;
    // Host resume
    `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    #20us;

    init_callback();
    bulk_in_xfer();
    bulk_out_xfer();
    #10us;
  endtask
endclass

class brt_usb_reset_handshake_quick_resume_vseq extends brt_usb_base_virtual_sequence;

  `brt_object_utils_begin(brt_usb_reset_handshake_quick_resume_vseq)
  `brt_object_utils_end

  function new(string name="brt_usb_reset_handshake_quick_resume_vseq");
    super.new(name);
  endfunction

  virtual task body();
    brt_usb_base_control_xfer_sequence              ctrl_seq;
    brt_usb_link_service_reset_sequence             reset_seq;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;
    brt_usb_agent_wait_for_link_usb_20_state_virtual_sequence wait_state;

    super.body();
    host_cfg.tdchbit = 2.5us;
    host_cfg.tdrsmdn = 1ms;
    dev_agt.cfg.tdrsmdn = 1ms;

    // Start
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::DEVICE_ATTACHED);
    // Reset device
    `brt_do_on(reset_seq, p_sequencer.link_service_sequencer) 

    `brt_info("DD", $sformatf("Wait for link state to ENABLE state"), UVM_LOW)
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    `brt_info("DD", $sformatf("link is ENABLE state"), UVM_LOW)

    #50us; 
    // reset 2nd time
    `brt_info("DD", $sformatf("link start to reset"), UVM_LOW)
    `brt_do_on(reset_seq, p_sequencer.link_service_sequencer) 
    `brt_info("DD", $sformatf("link is reseting"), UVM_LOW)
    // Wait ENABLE
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    `brt_info("DD", $sformatf("link is ENABLE state"), UVM_LOW)

    // let device enter suspend
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::SUSPENDED);

    #50us;
    // Host resume
    `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    #20us;

    init_callback();
    bulk_in_xfer();
    bulk_out_xfer();
    #10us;
  endtask
endclass

class brt_usb_dev_resume_vseq extends brt_usb_base_virtual_sequence;

  `brt_object_utils_begin(brt_usb_dev_resume_vseq)
  `brt_object_utils_end

  function new(string name="brt_usb_dev_resume_vseq");
    super.new(name);
  endfunction

  virtual task body();
    brt_usb_base_control_xfer_sequence              ctrl_seq;
    brt_usb_link_service_reset_sequence             reset_seq;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;
    brt_usb_agent_wait_for_link_usb_20_state_virtual_sequence wait_state;

    // Start
    super.body();

    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::DEVICE_ATTACHED);
    // Reset device
    `brt_do_on(reset_seq, p_sequencer.link_service_sequencer) 

    `brt_info("DD", $sformatf("Wait for link state to ENABLE state"), UVM_LOW)
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    `brt_info("DD", $sformatf("link is ENABLE state"), UVM_LOW)

    #50us; 
    // let device enter suspend
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::SUSPENDED);

    #50us;
    // dev resume
    `brt_do_on(resume_seq, dev_agt.link_service_sequencer) 
    wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);
    #20us;

    init_callback();
    bulk_in_xfer();
    bulk_out_xfer();
    #10us;
  endtask
endclass

// test mode
class brt_usb_testmode_nak_sequence extends brt_sequence #(brt_usb_packet);
    `brt_object_utils(brt_usb_testmode_nak_sequence)
    `brt_declare_p_sequencer (brt_usb_packet_sequencer)
    bit     terminate;
    bit     crc5_err;

    function new(string name="brt_usb_testmode_nak_sequence");
        super.new(name);
    endfunction

    virtual task body();
        forever begin
            req = brt_usb_packet::type_id::create();
            req.speed = brt_usb_types::FS;  // For randomize inter packet delay
            req.rx_to_tx = 0;         // For randomize inter packet delay
            start_item(req);
            if (!req.randomize() with {pid_name == brt_usb_packet::IN; func_address == 10; endp == 3;})
              `brt_fatal(get_name(), "randomize error")
            
            req.need_rsp = 1;  // Need data response
            // CRC5 err
            if (crc5_err) begin
                req.token_crc5 += $urandom_range(1,2**5-1);
                req.need_rsp = 0;  // Need data response
            end
            finish_item(req);
            get_response(rsp);
            if (req.need_rsp == 1) begin
                if (rsp.pid_format[3:0] == 4'ha) begin
                    `brt_info ("TESTMODE","Receive a NAK packet", UVM_LOW)
                end 
                else begin
                    `brt_error ("TESTMODE","Receive non-NAK packet")
                end
            end
            else begin
                #166666ps;
            end

            if (terminate) break;
        end
    endtask
endclass

class brt_usb_testmode_data0_sequence extends brt_sequence #(brt_usb_packet);
    `brt_object_utils(brt_usb_testmode_data0_sequence)
    `brt_declare_p_sequencer (brt_usb_packet_sequencer)
    bit     terminate;
    bit     crc5_err;

    function new(string name="brt_usb_testmode_data0_sequence");
        super.new(name);
    endfunction

    virtual task body();
        forever begin
            req = brt_usb_packet::type_id::create();
            req.speed = brt_usb_types::FS;  // For randomize inter packet delay
            req.rx_to_tx = 0;         // For randomize inter packet delay
            start_item(req);
            if (!req.randomize() with {pid_name == brt_usb_packet::IN; func_address == 10; endp == 3;})
              `brt_fatal(get_name(), "randomize error")
            
            req.need_rsp = 0;  // Need data response
            finish_item(req);
            get_response(rsp);
            #5us;

            if (terminate) break;
        end
    endtask
endclass

class brt_usb_testmode_nak_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_testmode_nak_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_testmode_nak_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1;
        host_cfg.remote_device_cfg[0].device_address = 10;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_testmode_nak_sequence   testmode_nak_seq;
        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        for (int i = 1; i < 1000; i++) begin
            dev_util_cb.add_inject_err (
                                          .addr          (  10                      ) // = 'hff
                                         ,.epnum         (  3                       ) // = 'h1f
                                         ,.dir           (  1                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       ( i                        ) // = 'b11
                                         );
        end
        
        testmode_nak_seq = new();
        mult_sb.dis_all = 1;
        fork
            begin
                testmode_nak_seq.start(p_sequencer.brt_usb_20_pkt_sequencer);
            end
            begin
                #100us;
                testmode_nak_seq.terminate = 1;
            end
        join
        
    endtask
endclass

class brt_usb_testmode_crc5err_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_testmode_crc5err_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_testmode_crc5err_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1;
        host_cfg.remote_device_cfg[0].device_address = 10;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_testmode_nak_sequence   testmode_nak_seq;
        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        for (int i = 1; i < 1000; i++) begin
            dev_util_cb.add_inject_err (
                                          .addr          (  10                      ) // = 'hff
                                         ,.epnum         (  3                       ) // = 'h1f
                                         ,.dir           (  1                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       ( i                        ) // = 'b11
                                         );
        end
        
        testmode_nak_seq = new();
        mult_sb.dis_all = 1;
        fork
            begin
                testmode_nak_seq.crc5_err = 1;
                testmode_nak_seq.start(p_sequencer.brt_usb_20_pkt_sequencer);
            end
            begin
                #10us;
                testmode_nak_seq.crc5_err = 0;
            end
            begin
                #100us;
                testmode_nak_seq.terminate = 1;
            end
        join
        
    endtask
endclass

class brt_usb_testmode_data0_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_testmode_data0_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_testmode_data0_vseq");
        super.new(name);
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1;
        host_cfg.remote_device_cfg[0].device_address = 10;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_testmode_data0_sequence   testmode_data0_seq;
        int                               num_data0;
        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0     ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        testmode_data0_seq = new();
        mult_sb.dis_all = 1;
        fork
            begin
                testmode_data0_seq.start(p_sequencer.brt_usb_20_pkt_sequencer);
            end
            fork
                forever begin
                    wait (p_sequencer.agt.prot.pkt_q.size() > 0);
                    if (p_sequencer.agt.prot.pkt_q[0].pid_format[3:0] == 4'h3) begin
                        `brt_info ("CHKP", "Receive a DATA0 packet in receiving channel", UVM_LOW) 
                        num_data0++;
                    end
                    else begin
                        `brt_error ("CHKP", "Receive a non-DATA0 packet in receiving channel") 
                    end
                    void'(p_sequencer.agt.prot.pkt_q.pop_front());
                end
            join_none
            begin
                #100us;
                testmode_data0_seq.terminate = 1;
            end
        join
        
        if (num_data0 < 10) begin
             `brt_error ("CHKP", "Not receive enough DATA0 packet in receiving channel") 
        end 
    endtask
endclass


// BULK zero length
class brt_usb_bulk_in_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_in_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_in_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            bulk_in_xfer (.set_ep_num(), .set_payload_size(0));
            #1us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            bulk_out_xfer (.set_ep_num(), .set_payload_size(0));
            #1us;
        end
    join
  endtask
endclass

// CONTROL SETUP

class brt_usb_control_2stage_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_2stage_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_2stage_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  0                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  0                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  0                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  0                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  0                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.pid_err       (  1                       ) // = 'b11
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_crc5err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_crc5err_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_crc5err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (  1                       ) // = 'b11
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (  1                       ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_deserr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_deserr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_deserr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  17                      ) // = 'hff
                                 ,.epnum         (  4                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = 'b11
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (                          ) // = 'hff
                                 ,.epnum         (                          ) // = 'h1f
                                 ,.dir           (                          ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (  17                      ) // = 'hff
                                         ,.new_epnum     (  4                       ) // = 'h1f
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = 'b11
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.new_pid       (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_eoperr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_eoperr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_eoperr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    dev_agt.link.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = 'b11
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.eop_length    ( host_cfg.speed == brt_usb_types::HS? 16:8                       ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_data0_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_data0_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_data0_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.pid_err       (  1                       ) // = 'b11
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_data0_crc16err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_data0_crc16err_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_data0_crc16err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc16_err     (  1                       ) // = 'b11
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (  1                       ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_data0_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_data0_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_data0_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_data0_bitstufferr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_data0_bitstufferr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_data0_bitstufferr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.bit_stuff_err (  1                       ) // = 'b11
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (  1                       ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_data0_eoperr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_data0_eoperr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_data0_eoperr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.eop_length    (  host_cfg.speed == brt_usb_types::HS? 16:8) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_data0_babbleerr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_data0_babbleerr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_data0_babbleerr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  9                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (  9                       ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.eop_length    (                          ) // = 'b11
                                         ,.rty           (  1                       ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_nak_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_nak_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_NAK"), .new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_nyet_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_nyet_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_nyet_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc16_err     (  1                       ) // = 'b11
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_stall_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_stall_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_STALL"), .new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("EP_HALT"), .new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         );

            mult_sb.disable_sb (0,0);                                         
            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_dev_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_dev_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_dev_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_STALL"), .new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("EP_HALT"), .new_severity(UVM_WARNING));

    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (  1                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

class brt_usb_control_setup_dev_eoperr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_setup_dev_eoperr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_setup_dev_eoperr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_data_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("p2d_seq"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.mon.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.mon.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.udriver.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_STALL"), .new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("EP_HALT"), .new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL), .id("x2p_seq0"), .new_severity(UVM_WARNING));

    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.eop_length    (  host_cfg.speed == brt_usb_types::HS ? 0 : 8) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(0));
        end
    join
  endtask
endclass

// 3 STAGE IN

class brt_usb_control_3stage_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_3stage_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_3stage_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_token_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_token_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_token_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_token_deserr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_token_deserr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_token_deserr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  17                      ) // = 'hff
                                 ,.epnum         (  4                       ) // = 'h1f
                                 ,.dir           (                          ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.new_addr      (  17                      ) // = 'hff
                                         ,.new_epnum     (  4                       ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  5                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_token_toggleerr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_token_toggleerr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_token_toggleerr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  5                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_data_nak_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_data_nak_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_data_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       ( 5                        ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_data_nyet_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_data_nyet_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_data_nyet_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       ( 5                        ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_data_stall_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_data_stall_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_data_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_STALL"), .new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("EP_HALT"), .new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       ( 5                        ) // = 'b11
                                         );
            mult_sb.disable_sb (0,0);                                         
            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_ack_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_ack_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_ack_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING x2p_seq0
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (  1                       ) // = -1
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          )
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.rty           (  1                       ) // = 'b11
                                         ,.pkt_idx       (  5                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_ack_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_ack_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_ack_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_IN_RSP"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  12                      ) // = -1
                                 ,.pkt_idx       (                          )
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (  12                      ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  5                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_in_ack_timeout_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_ack_timeout_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_ack_timeout_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_IN_RSP"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.pkt_idx       (  5                       ) // = 'b11
                                         );
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  5                       ) // = 'b11
                                         );

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.pkt_dly       (  50us                    ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(host_cfg.speed == brt_usb_types::LS ? 39:300));
        end
    join
  endtask
endclass

class brt_usb_control_in_littledata_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_littledata_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_littledata_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_IN_RSP"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (                          )
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            ctrl_xfer (.set_dir(1), .set_payload_size(300), .set_dev_payload_size(128));
        end
    join
  endtask
endclass

class brt_usb_control_in_alignwozero_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_alignwozero_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_alignwozero_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_IN_RSP"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 1;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            ctrl_xfer (.set_dir(1), .set_payload_size(128), .set_dev_payload_size(128));
        end
    join
  endtask
endclass

class brt_usb_control_in_alignwzero_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_alignwzero_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_alignwzero_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_IN_RSP"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            ctrl_xfer (.set_dir(1), .set_payload_size(128), .set_dev_payload_size(128));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_token_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_token_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_token_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (  1                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_token_deserr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_token_deserr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_token_deserr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  12                      ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (                          ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (                          ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.new_addr      (  12                      ) // = 'hff
                                         ,.new_epnum     (  1                       ) // = 'hff
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_token_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_token_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_token_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (                          ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (                          ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::IN      ) // = 'hff
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_data_crc16err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_data_crc16err_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_data_crc16err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.crc16_err     (  1                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (  1                       ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_data_babbleerr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_data_babbleerr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_data_babbleerr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1                       ) // = -1
                                 ,.crc16_err     (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            //chk_pkt.add_chk_pnt (
            //                      .addr          (  127                     ) // = 'hff
            //                     ,.epnum         (  0                       ) // = 'h1f
            //                     ,.dir           (  0                       ) // = 'b11
            //                     ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
            //                     ,.data_size     (                          ) // = -1
            //                     ,.pkt_idx       (  5                       ) // = -1
            //                     );
            //chk_pkt.add_chk_pnt (
            //                      .addr          (  127                     ) // = 'hff
            //                     ,.epnum         (  0                       ) // = 'h1f
            //                     ,.dir           (  0                       ) // = 'b11
            //                     ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
            //                     ,.data_size     (  0                       ) // = -1
            //                     ,.pkt_idx       (  5                       ) // = -1
            //                     );
            //chk_pkt.add_chk_pnt (
            //                      .addr          (  127                     ) // = 'hff
            //                     ,.epnum         (  0                       ) // = 'h1f
            //                     ,.dir           (  0                       ) // = 'b11
            //                     ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
            //                     ,.data_size     (                          ) // = -1
            //                     );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.data_size     (  1                       ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.rty           (                          ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(1), .set_payload_size(100));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_control_statusout_ack_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_ack_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_ack_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING   
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (  1                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  host_cfg.speed == brt_usb_types::LS ? 15 : 4 ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_ack_eoperr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_ack_eoperr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_ack_eoperr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING   
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_data_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("p2d_seq"),.new_severity(UVM_WARNING));
    dev_agt.mon.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.mon.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.udriver.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.eop_length    (  host_cfg.speed == brt_usb_types::HS? 0:8 ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_ack_nak_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_ack_nak_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_ack_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING   
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_ack_nyet_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_ack_nyet_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_ack_nyet_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING   
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_control_statusout_ack_stall_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_statusout_ack_stall_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_statusout_ack_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING   
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  4                       ) // = 'b11
                                         );
            mult_sb.disable_sb (0,0);                                         
            ctrl_xfer (.set_dir(1), .set_payload_size(100));
        end
    join
  endtask
endclass


class brt_usb_control_in_dev_data_errpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_dev_data_errpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_dev_data_errpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  ( 1                        ) // = 'b11
                                         ,.pkt_idx       ( 2                        ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(140));
        end
    join
  endtask
endclass

class brt_usb_control_in_dev_data_errcrc16_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_dev_data_errcrc16_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_dev_data_errcrc16_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (  1                       ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  ( 1                        ) // = 'b11
                                         ,.pkt_idx       ( 2                        ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(140));
        end
    join
  endtask
endclass

class brt_usb_control_in_dev_data_wrong_toggle_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_dev_data_wrong_toggle_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_dev_data_wrong_toggle_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.rty           ( 1                        ) // = 'b11
                                         ,.pkt_idx       ( 2                        ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(140));
        end
    join
  endtask
endclass

class brt_usb_control_in_dev_data_bitstuff_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_dev_data_bitstuff_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_dev_data_bitstuff_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_data_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("p2d_seq"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (  1                       ) // = 'b11
                                         ,.need_timeout  ( 1                        ) // = 'b11
                                         ,.pkt_idx       ( 2                        ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(140));
        end
    join
  endtask
endclass

class brt_usb_control_in_dev_data_erreop_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_dev_data_erreop_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_dev_data_erreop_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_data_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("p2d_seq"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    dev_agt.mon.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.mon.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.udriver.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.eop_length    (  host_cfg.speed == brt_usb_types::HS? 0:8 ) // = 'b11
                                         ,.need_timeout  ( 1                        ) // = 'b11
                                         ,.pkt_idx       ( 2                        ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(140));
        end
    join
  endtask
endclass

class brt_usb_control_in_dev_data_babble_errcrc16_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_in_dev_data_babble_errcrc16_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_in_dev_data_babble_errcrc16_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // Data stage
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (  1025                    ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (  1                       ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  ( 1                        ) // = 'b11
                                         ,.pkt_idx       ( 2                        ) // = 'b11
                                         );
            ctrl_xfer (.set_dir(1), .set_payload_size(140));
        end
    join
  endtask
endclass


// 3 STAGE OUT
class brt_usb_control_3stage_out_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_3stage_out_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_3stage_out_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );

            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_token_crc5err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_token_crc5err_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_token_crc5err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (  1                       ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (  1                       ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_token_deserr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_token_deserr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_token_deserr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  12                      ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (                          ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.new_addr      (  12                      ) // = 'hff
                                         ,.new_epnum     (  5                       ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_token_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_token_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_token_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_data_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_data_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_data_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_STALL"), .new_severity(UVM_WARNING));
    //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("EP_HALT"), .new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pid_err       (  1                       ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            //host_util_cb.add_inject_err (
            //                              .addr          (  127                     ) // = 'hff
            //                             ,.epnum         (  0                       ) // = 'h1f
            //                             ,.dir           (  0                       ) // = 'b11
            //                             ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
            //                             ,.new_pid       (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
            //                             ,.new_addr      (                          ) // = 'hff
            //                             ,.new_epnum     (                          ) // = 'h1f
            //                             ,.data_size     (                          ) // = -1
            //                             ,.pkt_err       (                          ) // = 'b00
            //                             ,.pid_err       (                          ) // = 'b11
            //                             ,.crc5_err      (                          ) // = 'b11
            //                             ,.crc16_err     (                          ) // = 'b11
            //                             ,.bit_stuff_err (                          ) // = 'b11
            //                             ,.need_timeout  (  1                       ) // = 'b11
            //                             ,.pkt_idx       (  3                       ) // = 'b11
            //                             );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_data_crc16err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_data_crc16err_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_data_crc16err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_STALL"), .new_severity(UVM_WARNING));
    //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("EP_HALT"), .new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.crc16_err     (  1                       ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            //host_util_cb.add_inject_err (
            //                              .addr          (  127                     ) // = 'hff
            //                             ,.epnum         (  0                       ) // = 'h1f
            //                             ,.dir           (  0                       ) // = 'b11
            //                             ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
            //                             ,.new_pid       (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
            //                             ,.new_addr      (                          ) // = 'hff
            //                             ,.new_epnum     (                          ) // = 'h1f
            //                             ,.data_size     (                          ) // = -1
            //                             ,.pkt_err       (                          ) // = 'b00
            //                             ,.pid_err       (                          ) // = 'b11
            //                             ,.crc5_err      (                          ) // = 'b11
            //                             ,.crc16_err     (                          ) // = 'b11
            //                             ,.bit_stuff_err (                          ) // = 'b11
            //                             ,.need_timeout  (  1                       ) // = 'b11
            //                             ,.pkt_idx       (  3                       ) // = 'b11
            //                             );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (  1                       ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_data_toggleerr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_data_toggleerr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_data_toggleerr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_STALL"), .new_severity(UVM_WARNING));
    //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("EP_HALT"), .new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.crc16_err     (                          ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            //host_util_cb.add_inject_err (
            //                              .addr          (  127                     ) // = 'hff
            //                             ,.epnum         (  0                       ) // = 'h1f
            //                             ,.dir           (  0                       ) // = 'b11
            //                             ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
            //                             ,.new_pid       (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
            //                             ,.new_addr      (                          ) // = 'hff
            //                             ,.new_epnum     (                          ) // = 'h1f
            //                             ,.data_size     (                          ) // = -1
            //                             ,.pkt_err       (                          ) // = 'b00
            //                             ,.pid_err       (                          ) // = 'b11
            //                             ,.crc5_err      (                          ) // = 'b11
            //                             ,.crc16_err     (                          ) // = 'b11
            //                             ,.bit_stuff_err (                          ) // = 'b11
            //                             ,.need_timeout  (  1                       ) // = 'b11
            //                             ,.pkt_idx       (  3                       ) // = 'b11
            //                             );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_data_bistufferr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_data_bistufferr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_data_bistufferr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.bit_stuff_err (  1                       ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            //host_util_cb.add_inject_err (
            //                              .addr          (  127                     ) // = 'hff
            //                             ,.epnum         (  0                       ) // = 'h1f
            //                             ,.dir           (  0                       ) // = 'b11
            //                             ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
            //                             ,.new_pid       (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
            //                             ,.new_addr      (                          ) // = 'hff
            //                             ,.new_epnum     (                          ) // = 'h1f
            //                             ,.data_size     (                          ) // = -1
            //                             ,.pkt_err       (                          ) // = 'b00
            //                             ,.pid_err       (                          ) // = 'b11
            //                             ,.crc5_err      (                          ) // = 'b11
            //                             ,.crc16_err     (                          ) // = 'b11
            //                             ,.bit_stuff_err (                          ) // = 'b11
            //                             ,.need_timeout  (  1                       ) // = 'b11
            //                             ,.pkt_idx       (  3                       ) // = 'b11
            //                             );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (  1                       ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_data_babbleerr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_data_babbleerr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_data_babbleerr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  1025                    ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            //host_util_cb.add_inject_err (
            //                              .addr          (  127                     ) // = 'hff
            //                             ,.epnum         (  0                       ) // = 'h1f
            //                             ,.dir           (  0                       ) // = 'b11
            //                             ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
            //                             ,.new_pid       (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
            //                             ,.new_addr      (                          ) // = 'hff
            //                             ,.new_epnum     (                          ) // = 'h1f
            //                             ,.data_size     (                          ) // = -1
            //                             ,.pkt_err       (                          ) // = 'b00
            //                             ,.pid_err       (                          ) // = 'b11
            //                             ,.crc5_err      (                          ) // = 'b11
            //                             ,.crc16_err     (                          ) // = 'b11
            //                             ,.bit_stuff_err (                          ) // = 'b11
            //                             ,.need_timeout  (  1                       ) // = 'b11
            //                             ,.pkt_idx       (  3                       ) // = 'b11
            //                             );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (  1025                    ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_dev_ack_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_dev_ack_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_dev_ack_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pid_err       (  1                       ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (  1                       ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_dev_ack_eoperr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_dev_ack_eoperr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_dev_ack_eoperr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_data_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("p2d_seq"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.mon.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.mon.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    host_agt.udriver.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (  1                       ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.eop_length    (  host_cfg.speed == brt_usb_types::HS? 0:8 ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_dev_nak_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_dev_nak_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_dev_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_dev_nyet_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_dev_nyet_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_dev_nyet_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  8                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_dev_stall_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_dev_stall_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_dev_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("RCV_STALL"), .new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR), .id("EP_HALT"), .new_severity(UVM_WARNING));

    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.new_addr      (                          ) // = 'hff
                                         ,.new_epnum     (                          ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = 'b11
                                         );

            mult_sb.disable_sb (0,0);                                         
            ctrl_xfer (.set_dir(0), .set_payload_size(300));
        end
    join
  endtask
endclass

class brt_usb_control_out_allignwozero_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_allignwozero_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_allignwozero_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 1;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_out_allignwzero_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_out_allignwzero_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_out_allignwzero_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_token_crc5err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_token_crc5err_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_token_crc5err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (  1                       ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (  1                       ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_token_deserr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_token_deserr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_token_deserr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq1"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq1"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  12                      ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (                          ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.new_addr      (  12                      ) // = 'h1f
                                         ,.new_epnum     (  1                       ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_token_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_token_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_token_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::OUT     ) // = 'h1f
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_data_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_data_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_data_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // disable monitor checker
    host_cfg.ignore_mon_host_err = 1;
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (  1                       ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_data_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_data_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_data_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.rty           (  1                       ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_data_babbleerr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_data_babbleerr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_data_babbleerr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1                       ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.data_size     (  1                       ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_data_nak_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_data_nak_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_data_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_data_stall_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_data_stall_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_data_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            mult_sb.disable_sb (0,0);                                         
            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_ack_piderr_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_ack_piderr_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_ack_piderr_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pid_err       (  1                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.crc5_err      (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (                          ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

class brt_usb_control_status_ack_wrongpid_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_status_ack_wrongpid_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_control_status_ack_wrongpid_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change ERROR to WARNING
    host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq0"),.new_severity(UVM_WARNING));
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_IN_RSP"),.new_severity(UVM_WARNING));
    //dev_agt.link.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("brt_usb_link"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //host_agt.ulayer.link_mon.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("link_mon"),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
    // Change config
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[0].allow_aligned_transfer_without_zero_length = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
        
                         ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // zero length
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 );
            // Status
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  6                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.crc5_err      (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                       ) // = -1
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (  7                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.crc5_err      (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  0                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  6                       ) // = 'b11
                                         );

            ctrl_xfer (.set_dir(0), .set_payload_size(64*3));
        end
    join
  endtask
endclass

// CONTROL random
class brt_usb_control_random_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_control_random_vseq)
  `uvm_object_utils_end
  rand int  mps;
  rand int  xfer_size;
  constraint reasonable_mps {
      mps inside {8, 64};
  };
  constraint reasonable_xfer_size {
      xfer_size dist {0 := 1, [1:300] :/ 2};
  };

  function new(string name="brt_usb_control_random_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    // Change config
    host_cfg.remote_device_cfg[0].device_address = $urandom_range (0,127);
    dev_addr = host_cfg.remote_device_cfg[0].device_address;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            chk_pkt.add_chk_pnt (
                                  .addr          (  dev_addr                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::SETUP   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  dev_addr                     ) // = 'hff
                                 ,.epnum         (  0                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            repeat (16) begin
                this.randomize();
                host_cfg.remote_device_cfg[0].endpoint_cfg[0].max_packet_size = mps;
                #1;
                ctrl_xfer (.set_dir(), .set_payload_size(xfer_size));
            end
        end
    join
  endtask
endclass



// BULK IN
class brt_usb_bulk_in_mps8_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_in_mps8_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_in_mps8_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = 8;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_in_xfer (.set_payload_size(1500));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_mps64_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_in_mps64_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_in_mps64_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = 64;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_in_xfer (.set_payload_size(1499));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_mps512_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_in_mps512_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_in_mps512_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = 512;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  512                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_in_xfer (.set_payload_size(1499));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_mps1024_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_in_mps1024_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_in_mps1024_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_in_xfer (.set_payload_size(2499));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_align_short_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_in_align_short_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_in_align_short_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                        ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_in_xfer (.set_payload_size(3*1024),.set_dev_payload_size(1*1024));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_align_wo_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_in_align_wo_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_in_align_wo_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 1;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_in_xfer (.set_payload_size(3*1024),.set_dev_payload_size(3*1024));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_align_w_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_in_align_w_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_in_align_w_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                        ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_in_xfer (.set_payload_size(1*1024),.set_dev_payload_size(1*1024));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_token_pid_err_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_bulk_in_token_pid_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_in_token_pid_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  $urandom_range(1,3)     ) // = 'b11
                                         );


            repeat (3)
                bulk_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_token_crc5_err_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_bulk_in_token_crc5_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_in_token_crc5_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (  1                       ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  $urandom_range(1,3)     ) // = 'b11
                                         );


            repeat (3)
                bulk_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_token_rty_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_bulk_in_token_rty_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_in_token_rty_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    dev_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    host_agt.clear_ep_toggle (.epnum(1), .dir(1));
    dev_agt.clear_ep_toggle (.epnum(1), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            repeat (3)
                bulk_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_token_dev_timeout_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_bulk_in_token_dev_timeout_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_in_token_dev_timeout_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    dev_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    host_agt.clear_ep_toggle (.epnum(1), .dir(1));
    dev_agt.clear_ep_toggle (.epnum(1), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.drop          (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            repeat (3)
                bulk_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_token_dev_pid_err_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_bulk_in_token_dev_pid_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_in_token_dev_pid_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    dev_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    host_agt.clear_ep_toggle (.epnum(1), .dir(1));
    dev_agt.clear_ep_toggle (.epnum(1), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.drop          (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            repeat (3)
                bulk_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_nak_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_bulk_in_nak_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_in_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (                          ) // = 'b11
                                         );

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (                          ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (                          ) // = 'b11
                                         );

            repeat (1)
                bulk_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_bulk_in_stall_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_bulk_in_stall_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_in_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[1].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(1), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  1                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (                          ) // = 'b11
                                         );

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  1                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (                          ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (                          ) // = 'b11
                                         );
            mult_sb.dis_all = 1;
            bulk_in_xfer (.set_payload_size(xfer_size));
            host_agt.clear_halt_status(.epnum(1), .dir(1));
            dev_agt.abort_transfer(.epnum(1), .dir(1));
            mult_sb.dis_all = 0;
            bulk_in_xfer (.set_payload_size(xfer_size));
            //dev_agt.clear_halt_status(.epnum(1), .dir(1));
        end
    join
  endtask
endclass

// BULK OUT
class brt_usb_bulk_out_mps8_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_mps8_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_mps8_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = 8;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_out_xfer (.set_payload_size(500));
            bulk_out_xfer (.set_payload_size(1500));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_mps64_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_mps64_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_mps64_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = 64;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_out_xfer (.set_payload_size(499));
            bulk_out_xfer (.set_payload_size(1499));
        end
    join
  endtask
endclass

class brt_usb_bulk_out_mps512_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_mps512_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_mps512_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = 512;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  512                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_out_xfer (.set_payload_size(1499));
        end
    join
  endtask
endclass

class brt_usb_bulk_out_mps1024_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_mps1024_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_mps1024_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_out_xfer (.set_payload_size(2499));
        end
    join
  endtask
endclass

class brt_usb_bulk_out_align_wo_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_align_wo_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_align_wo_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 1;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_out_xfer (.set_payload_size(3*1024),.set_dev_payload_size(3*1024));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_align_w_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_align_w_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_align_w_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                        ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            bulk_out_xfer (.set_payload_size(1*1024),.set_dev_payload_size(1*1024));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_nyet_w_ping_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_nyet_w_ping_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_nyet_w_ping_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::PING    ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = -1
                                         );

            bulk_out_xfer (.set_payload_size(5*1024),.set_dev_payload_size(5*1024));
        end
    join
  endtask
endclass

class brt_usb_bulk_out_nyet_wo_ping_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_nyet_wo_ping_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_bulk_out_nyet_wo_ping_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = 1024;
    host_cfg.ping_support = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                    ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                    ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = -1
                                         );

            bulk_out_xfer (.set_payload_size(5*1024),.set_dev_payload_size(5*1024));
        end
    join
  endtask
endclass

class brt_usb_bulk_out_pid_err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_pid_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_out_pid_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(2), .dir(0));
    host_agt.clear_ep_toggle (.epnum(2), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(2), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.pid_err       (  1                       ) // = -1
                                 ,.pkt_idx       (  1                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  idx%2?brt_usb_packet::DATA0:brt_usb_packet::DATA1 ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (3)
                bulk_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_crc5_err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_crc5_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_out_crc5_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(2), .dir(0));
    host_agt.clear_ep_toggle (.epnum(2), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(2), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (  1                       ) // = -1
                                 ,.pkt_idx       (  1                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (  1                       ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  idx%2?brt_usb_packet::DATA0:brt_usb_packet::DATA1 ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (3)
                bulk_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_crc16_err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_crc16_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_out_crc16_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(2), .dir(0));
    host_agt.clear_ep_toggle (.epnum(2), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(2), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (                          ) // = brt_usb_packet::EXT
                                 ,.crc16_err     (  1                       ) // = -1
                                 ,.pkt_idx       (  1                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  idx%2?brt_usb_packet::DATA0:brt_usb_packet::DATA1 ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (  1                       ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (3)
                bulk_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_timeout_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_timeout_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_out_timeout_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(2), .dir(0));
    host_agt.clear_ep_toggle (.epnum(2), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(2), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  idx%2?brt_usb_packet::DATA0:brt_usb_packet::DATA1 ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (3)
                bulk_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_nak_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_nak_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_out_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = mps;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_num_nak_per_transfer = 1000;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(2), .dir(0));
    dev_util_cb.reset_index (.addr(127), .epnum(2), .dir(0));
    host_agt.clear_ep_toggle (.epnum(2), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(2), .dir(0));
    xfer_size = 1000;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            for(int i = 0; i<1000;i++)
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  i                       ) // = 'b11
                                         );

            fork begin
                #500us;
                host_agt.ulayer.x2p_seq[2].xfer_terminated = 1;
            end join_none

            repeat (1)
                bulk_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_bulk_out_stall_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_bulk_out_stall_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {8, 64, 128, 256, 512, 1024};
  };

  function new(string name="brt_usb_bulk_out_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[2].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(2), .dir(0));
    dev_util_cb.reset_index (.addr(127), .epnum(2), .dir(0));
    host_agt.clear_ep_toggle (.epnum(2), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(2), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  2                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  2                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            mult_sb.dis_all = 1;
            repeat (1) begin
                bulk_out_xfer (.set_payload_size(xfer_size));
            end
            host_agt.clear_halt_status(.epnum(2), .dir(0));
            #10us;
        end
    join
  endtask
endclass

// INTERRUPT IN
class brt_usb_int_in_mps8_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_mps8_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_mps8_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 8;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(100));
        end
    join
  endtask
endclass

class brt_usb_int_in_mps64_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_mps64_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_mps64_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 64;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(499));
        end
    join
  endtask
endclass

class brt_usb_int_in_mps512_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_mps512_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_mps512_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 512;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  512                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(1499));
        end
    join
  endtask
endclass

class brt_usb_int_in_mps1024_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_mps1024_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_mps1024_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 1024;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_burst_size = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(2499));
        end
    join
  endtask
endclass

class brt_usb_int_in_mps1024_burst1_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_mps1024_burst1_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_mps1024_burst1_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 1024;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_burst_size = 1;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(2499));
        end
    join
  endtask
endclass

class brt_usb_int_in_mps1024_burst2_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_mps1024_burst2_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_mps1024_burst2_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 1024;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_burst_size = 2;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(2499));
        end
    join
  endtask
endclass

class brt_usb_int_in_align_short_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_align_short_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_align_short_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                        ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(3*1024),.set_dev_payload_size(1*1024));
        end
    join
  endtask
endclass

class brt_usb_int_in_align_wo_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_align_wo_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_align_wo_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 1;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(3*1024),.set_dev_payload_size(3*1024));
        end
    join
  endtask
endclass

class brt_usb_int_in_align_w_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_in_align_w_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_in_align_w_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                        ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_in_xfer (.set_payload_size(1*1024),.set_dev_payload_size(1*1024));
        end
    join
  endtask
endclass

class brt_usb_int_in_token_pid_err_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_int_in_token_pid_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_in_token_pid_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(5), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  5                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  $urandom_range(1,2)     ) // = 'b11
                                         );


            repeat (2)
                interrupt_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_int_in_token_crc5_err_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_int_in_token_crc5_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_in_token_crc5_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(5), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  5                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (  1                       ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  $urandom_range(1,2)     ) // = 'b11
                                         );


            repeat (2)
                interrupt_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_int_in_token_rty_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_int_in_token_rty_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_in_token_rty_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(5), .dir(1));
    dev_util_cb.reset_index (.addr(127), .epnum(5), .dir(1));
    host_agt.clear_ep_toggle (.epnum(5), .dir(1));
    dev_agt.clear_ep_toggle (.epnum(5), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  5                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  5                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  1                       ) // = 'b11
                                         );

            repeat (1)
                interrupt_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_int_in_nak_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_int_in_nak_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_in_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(5), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  5                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (                          ) // = 'b11
                                         );

            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  5                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (                          ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (                          ) // = 'b11
                                         );

            repeat (1)
                interrupt_in_xfer (.set_payload_size(xfer_size));
        end
    join
  endtask
endclass

class brt_usb_int_in_stall_vseq extends brt_usb_base_virtual_sequence;
  `uvm_object_utils_begin(brt_usb_int_in_stall_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_in_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[5].max_packet_size = mps;
    reset_dev();

    xfer_size = host_cfg.speed == brt_usb_types::HS? 3333:555;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(5), .dir(1));
    xfer_size = 0;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  5                       ) // = 'h1f
                                 ,.dir           (  1                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  5                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (                          ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (                          ) // = 'b11
                                         );
            mult_sb.dis_all = 1;
            repeat (1)
                interrupt_in_xfer (.set_payload_size(xfer_size));

            host_agt.clear_halt_status(.epnum(5), .dir(1));
            //dev_agt.clear_halt_status(.epnum(5), .dir(1));
        end
    join
  endtask
endclass


// INTERRUPT OUT
class brt_usb_int_out_mps8_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_mps8_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_mps8_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 8;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  8                       ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_out_xfer (.set_payload_size(100));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_int_out_mps64_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_mps64_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_mps64_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 64;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  64                      ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_out_xfer (.set_payload_size(499));
        end
    join
  endtask
endclass

class brt_usb_int_out_mps512_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_mps512_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_mps512_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 512;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  512                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_out_xfer (.set_payload_size(1499));
        end
    join
  endtask
endclass

class brt_usb_int_out_mps1024_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_mps1024_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_mps1024_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 1024;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_burst_size  = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_out_xfer (.set_payload_size(2499));
        end
    join
  endtask
endclass

class brt_usb_int_out_mps1024_burst1_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_mps1024_burst1_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_mps1024_burst1_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 1024;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_burst_size  = 1;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_out_xfer (.set_payload_size(2499));
        end
    join
  endtask
endclass

class brt_usb_int_out_mps1024_burst2_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_mps1024_burst2_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_mps1024_burst2_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 1024;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_burst_size  = 2;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_out_xfer (.set_payload_size(2499));
        end
    join
  endtask
endclass

class brt_usb_int_out_align_wo_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_align_wo_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_align_wo_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 1;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_out_xfer (.set_payload_size(3*1024),.set_dev_payload_size(3*1024));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_int_out_align_w_zerolen_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_align_w_zerolen_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_align_w_zerolen_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  0                        ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);

            interrupt_out_xfer (.set_payload_size(1*1024),.set_dev_payload_size(1*1024));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_int_out_nyet_w_ping_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_nyet_w_ping_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_nyet_w_ping_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 1024;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::PING    ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  5                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = -1
                                         );

            interrupt_out_xfer (.set_payload_size(5*1024),.set_dev_payload_size(5*1024));
        end
    join
  endtask
endclass

class brt_usb_int_out_nyet_wo_ping_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_nyet_wo_ping_vseq)
  `uvm_object_utils_end

  function new(string name="brt_usb_int_out_nyet_wo_ping_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = 1024;
    host_cfg.ping_support = 0;
    reset_dev();
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                     ) // = -1
                                 ,.pkt_idx       (  2                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                    ) // = -1
                                 ,.pkt_idx       (  3                       ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                 ,.data_size     (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                 ,.data_size     (  1024                    ) // = -1
                                 ,.pkt_idx       (  4                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (  0                       ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  3                       ) // = -1
                                         );

            interrupt_out_xfer (.set_payload_size(5*1024),.set_dev_payload_size(5*1024));
        end
    join
  endtask
endclass

class brt_usb_int_out_pid_err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_pid_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_out_pid_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(6), .dir(0));
    host_agt.clear_ep_toggle (.epnum(6), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(6), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.pid_err       (  1                       ) // = -1
                                 ,.pkt_idx       (  1                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (  1                       ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  idx%2?brt_usb_packet::DATA0:brt_usb_packet::DATA1 ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (3)
                interrupt_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_int_out_crc5_err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_crc5_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_out_crc5_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(6), .dir(0));
    host_agt.clear_ep_toggle (.epnum(6), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(6), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::OUT      ) // = brt_usb_packet::EXT
                                 ,.crc5_err      (  1                       ) // = -1
                                 ,.pkt_idx       (  1                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (  1                       ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  idx%2?brt_usb_packet::DATA0:brt_usb_packet::DATA1 ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (3)
                interrupt_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_int_out_crc16_err_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_crc16_err_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_out_crc16_err_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(6), .dir(0));
    host_agt.clear_ep_toggle (.epnum(6), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(6), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (                          ) // = brt_usb_packet::EXT
                                 ,.crc16_err     (  1                       ) // = -1
                                 ,.pkt_idx       (  1                       ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  idx%2?brt_usb_packet::DATA0:brt_usb_packet::DATA1 ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (  1                       ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (3)
                interrupt_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_int_out_timeout_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_timeout_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_out_timeout_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(6), .dir(0));
    host_agt.clear_ep_toggle (.epnum(6), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(6), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // error injection
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );
            host_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  idx%2?brt_usb_packet::DATA0:brt_usb_packet::DATA1 ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.drop          (  1                       ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (3)
                interrupt_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_int_out_nak_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_nak_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_out_nak_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = mps;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(6), .dir(0));
    dev_util_cb.reset_index (.addr(127), .epnum(6), .dir(0));
    host_agt.clear_ep_toggle (.epnum(6), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(6), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::NAK     ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            repeat (2)
                interrupt_out_xfer (.set_payload_size(xfer_size));
            #10us;
        end
    join
  endtask
endclass

class brt_usb_int_out_stall_vseq extends brt_usb_base_virtual_sequence;

  `uvm_object_utils_begin(brt_usb_int_out_stall_vseq)
  `uvm_object_utils_end

  rand int  mps;
  int       xfer_size;
  int       idx;
  constraint reasonable_mps {
      mps inside {256, 512, 1024};
  };

  function new(string name="brt_usb_int_out_stall_vseq");
    super.new(name);
  endfunction

  virtual task body();
    super.body();
    this.randomize();
    host_cfg.remote_device_cfg[0].device_address = 127;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].allow_aligned_transfer_without_zero_length = 0;
    host_cfg.remote_device_cfg[0].endpoint_cfg[6].max_packet_size = mps;
    host_cfg.run = 0;
    #25ms;
    host_cfg.run = 1;
    reset_dev();
    xfer_size = host_cfg.speed == brt_usb_types::HS? $urandom_range (3000,5000):$urandom_range (300,500) ;
    idx = 2;
    start_xfer();
    host_util_cb.reset_index (.addr(127), .epnum(6), .dir(0));
    dev_util_cb.reset_index (.addr(127), .epnum(6), .dir(0));
    host_agt.clear_ep_toggle (.epnum(6), .dir(0));
    dev_agt.clear_ep_toggle (.epnum(6), .dir(0));
    xfer_size = 0;
    idx = 1;
    start_xfer();
  endtask

  virtual task start_xfer();
    brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

    // Start SOF
    `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
    `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
    `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)


    fork
        // CTRL
        begin
            // Checker
            chk_pkt = new("chk_pkt", host_util_cb);
            // data
            chk_pkt.add_chk_pnt (
                                  .addr          (  127                     ) // = 'hff
                                 ,.epnum         (  6                       ) // = 'h1f
                                 ,.dir           (  0                       ) // = 'b11
                                 ,.pid           (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                 ,.pid_err       (                          ) // = -1
                                 ,.pkt_idx       (                          ) // = -1
                                 );
            host_util_cb.add_chk_pkt(chk_pkt);
            // error injection
            dev_util_cb.add_inject_err (
                                          .addr          (  127                     ) // = 'hff
                                         ,.epnum         (  6                       ) // = 'h1f
                                         ,.dir           (                          ) // = 'b11
                                         ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                         ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                         ,.data_size     (                          ) // = -1
                                         ,.pkt_err       (                          ) // = 'b00
                                         ,.pid_err       (                          ) // = 'b11
                                         ,.crc5_err      (                          ) // = 'b11
                                         ,.crc16_err     (                          ) // = 'b11
                                         ,.bit_stuff_err (                          ) // = 'b11
                                         ,.need_timeout  (                          ) // = 'b11
                                         ,.pkt_idx       (  idx                     ) // = 'b11
                                         );

            mult_sb.dis_all = 1;
            repeat (1) begin
                interrupt_out_xfer (.set_payload_size(xfer_size));
            end
            host_agt.clear_halt_status(.epnum(6), .dir(0));
            #10us;
        end
    join
  endtask
endclass


// ISO IN
class brt_usb_iso_in_mps1_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_mps1_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_mps1_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(1));
        isochronous_in_xfer(.set_payload_size(1));
        isochronous_in_xfer(.set_payload_size(0));
        isochronous_in_xfer(.set_payload_size(0));
    endtask
endclass

class brt_usb_iso_in_mps8_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_mps8_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_mps8_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 8;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 8;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  8                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  8                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(8));
        isochronous_in_xfer(.set_payload_size(8));
        isochronous_in_xfer(.set_payload_size(0));
        isochronous_in_xfer(.set_payload_size(0));
    endtask
endclass

class brt_usb_iso_in_mps77_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_mps77_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_mps77_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 77;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 77;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  77                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  77                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(77));
        isochronous_in_xfer(.set_payload_size(77));
        isochronous_in_xfer(.set_payload_size(55));
        isochronous_in_xfer(.set_payload_size(55));
    endtask
endclass

class brt_usb_iso_in_mps512_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_mps512_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_mps512_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 512;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 512;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  512                     ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  512                     ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(512));
        isochronous_in_xfer(.set_payload_size(512));
        isochronous_in_xfer(.set_payload_size(0));
        isochronous_in_xfer(.set_payload_size(0));
    endtask
endclass

class brt_usb_iso_in_mps567_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_mps567_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_mps567_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 567;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 567;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  567                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  567                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(567));
        isochronous_in_xfer(.set_payload_size(567));
        isochronous_in_xfer(.set_payload_size(55));
        isochronous_in_xfer(.set_payload_size(55));
    endtask
endclass

class brt_usb_iso_in_mps1024_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_mps1024_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_mps1024_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(1024));
        isochronous_in_xfer(.set_payload_size(1024));
        isochronous_in_xfer(.set_payload_size(55));
        isochronous_in_xfer(.set_payload_size(55));
    endtask
endclass

class brt_usb_iso_in_burst2_mps513_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_burst2_mps513_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_burst2_mps513_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 513;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 513;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  513                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  513                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(1000));
        isochronous_in_xfer(.set_payload_size(1000));
    endtask
endclass

class brt_usb_iso_in_burst2_mps1024_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_burst2_mps1024_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_burst2_mps1024_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(1000));
        isochronous_in_xfer(.set_payload_size(2000));
    endtask
endclass

class brt_usb_iso_in_burst3_mps683_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_burst3_mps683_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_burst3_mps683_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 683;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 683;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  683                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  683                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  683                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  683                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(1700));
        isochronous_in_xfer(.set_payload_size(1700));
    endtask
endclass

class brt_usb_iso_in_burst3_mps1024_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_burst3_mps1024_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_burst3_mps1024_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(700));
        isochronous_in_xfer(.set_payload_size(1700));
        isochronous_in_xfer(.set_payload_size(2700));
    endtask
endclass

class brt_usb_iso_in_burst3_mps1024_token_pid_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_burst3_mps1024_token_pid_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_burst3_mps1024_token_pid_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  3                       ) // = 'h1f
                                     ,.dir           (  1                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (  1                       ) // = 'b11
                                     ,.crc5_err      (                          ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(2700));
        mult_sb.enable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(2700));
    endtask
endclass

class brt_usb_iso_in_burst3_mps1024_token_crc5_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_burst3_mps1024_token_crc5_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_burst3_mps1024_token_crc5_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  3                       ) // = 'h1f
                                     ,.dir           (  1                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (  1                       ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(2700));
        mult_sb.enable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(2700));
    endtask
endclass

class brt_usb_iso_in_burst3_mps1024_data_wrongpid_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_burst3_mps1024_data_wrongpid_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_burst3_mps1024_data_wrongpid_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        // Change ERROR to WARNING
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        dev_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  3                       ) // = 'h1f
                                     ,.dir           (  1                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                                     ,.new_pid       (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (                          ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (                          ) // = 'b11
                                     );
        
        mult_sb.disable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(2700));
        mult_sb.enable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(2700));
    endtask
endclass

class brt_usb_iso_in_burst3_mps1024_xfer_babble_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_burst3_mps1024_xfer_babble_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_burst3_mps1024_xfer_babble_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        // Change ERROR to WARNING x2p_seq3
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("x2p_seq3"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1000                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        dev_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  3                       ) // = 'h1f
                                     ,.dir           (  1                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                                     ,.data_size     (  1000                    ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (                          ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (                          ) // = 'b11
                                     );
        
        mult_sb.disable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(2700));
        mult_sb.enable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(2700));
    endtask
endclass

class brt_usb_iso_in_mps512_token_crc5_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_mps512_token_crc5_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_mps512_token_crc5_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 512;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 512;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  3                       ) // = 'h1f
                                     ,.dir           (  1                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (  1                       ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(500));
        mult_sb.enable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(500));
    endtask
endclass

class brt_usb_iso_in_mps512_token_pid_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_in_mps512_token_pid_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_mps512_token_pid_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 512;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 512;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  3                       ) // = 'h1f
                                     ,.dir           (  1                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::IN      ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (  1                       ) // = 'b11
                                     ,.crc5_err      (                          ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(500));
        mult_sb.enable_sb (3,1);                                         
        isochronous_in_xfer(.set_payload_size(500));
    endtask
endclass

// ISO OUT
class brt_usb_iso_out_mps1_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_mps1_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_mps1_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(1));
        isochronous_out_xfer(.set_payload_size(1));
        isochronous_out_xfer(.set_payload_size(0));
        isochronous_out_xfer(.set_payload_size(0));
        #1us;
    endtask
endclass

class brt_usb_iso_out_mps8_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_mps8_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_mps8_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 8;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 8;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  8                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  8                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(8));
        isochronous_out_xfer(.set_payload_size(8));
        isochronous_out_xfer(.set_payload_size(0));
        isochronous_out_xfer(.set_payload_size(0));
        #1us;
    endtask
endclass

class brt_usb_iso_out_mps77_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_mps77_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_mps77_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 77;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 77;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  77                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  77                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(77));
        isochronous_out_xfer(.set_payload_size(77));
        isochronous_out_xfer(.set_payload_size(55));
        isochronous_out_xfer(.set_payload_size(55));
        #1us;
    endtask
endclass

class brt_usb_iso_out_mps512_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_mps512_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_mps512_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 512;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 512;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  512                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  512                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  0                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(512));
        isochronous_out_xfer(.set_payload_size(512));
        isochronous_out_xfer(.set_payload_size(0));
        isochronous_out_xfer(.set_payload_size(0));
        #1us;
    endtask
endclass

class brt_usb_iso_out_mps567_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_mps567_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_mps567_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 567;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 567;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  567                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  567                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(567));
        isochronous_out_xfer(.set_payload_size(567));
        isochronous_out_xfer(.set_payload_size(55));
        isochronous_out_xfer(.set_payload_size(55));
        #1us;
    endtask
endclass

class brt_usb_iso_out_mps1024_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_mps1024_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_mps1024_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(1024));
        isochronous_out_xfer(.set_payload_size(1024));
        isochronous_out_xfer(.set_payload_size(55));
        isochronous_out_xfer(.set_payload_size(55));
        #1us;
    endtask
endclass

class brt_usb_iso_out_burst2_mps513_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_burst2_mps513_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_burst2_mps513_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 513;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 513;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  513                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  513                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(1000));
        isochronous_out_xfer(.set_payload_size(1000));
        #1us;
    endtask
endclass

class brt_usb_iso_out_burst2_mps1024_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_burst2_mps1024_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_burst2_mps1024_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 1;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA1   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(1000));
        isochronous_out_xfer(.set_payload_size(2000));
        #1us;
    endtask
endclass

class brt_usb_iso_out_burst3_mps683_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_burst3_mps683_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_burst3_mps683_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 683;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 683;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  683                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  683                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  683                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  683                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(1700));
        isochronous_out_xfer(.set_payload_size(1700));
        #1us;
    endtask
endclass

class brt_usb_iso_out_burst3_mps1024_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_burst3_mps1024_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_burst3_mps1024_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_out_xfer(.set_payload_size(2700));
        isochronous_out_xfer(.set_payload_size(2700));
        #1us;
    endtask
endclass

class brt_usb_iso_out_burst3_mps1024_token_pid_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_burst3_mps1024_token_pid_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_burst3_mps1024_token_pid_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  4                       ) // = 'h1f
                                     ,.dir           (  0                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (  1                       ) // = 'b11
                                     ,.crc5_err      (                          ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(2700));
        //mult_sb.enable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(2700));
        #1us;
    endtask
endclass

class brt_usb_iso_out_burst3_mps1024_token_crc5_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_burst3_mps1024_token_crc5_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_burst3_mps1024_token_crc5_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  4                       ) // = 'h1f
                                     ,.dir           (  0                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (  1                       ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(2700));
        //mult_sb.enable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(2700));
        #1us;
    endtask
endclass

class brt_usb_iso_out_burst3_mps1024_data_wrongpid_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_burst3_mps1024_data_wrongpid_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_burst3_mps1024_data_wrongpid_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        // Change ERROR to WARNING
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("d_x2p_seq4"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  4                       ) // = 'h1f
                                     ,.dir           (  0                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                                     ,.new_pid       (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (                          ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(2700));
        #1us;
        //mult_sb.enable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(2700));
        #1us;
    endtask
endclass

class brt_usb_iso_out_burst3_mps1024_xfer_babble_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_burst3_mps1024_xfer_babble_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_burst3_mps1024_xfer_babble_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        // Change ERROR to WARNING
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 2;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1000                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::MDATA   ) // = brt_usb_packet::EXT
                             ,.data_size     (  1024                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  4                       ) // = 'h1f
                                     ,.dir           (  0                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA2   ) // = brt_usb_packet::EXT
                                     ,.data_size     (  1000                    ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (                          ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (                          ) // = 'b11
                                     );
        
        mult_sb.disable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(2700));
        #1us;
        mult_sb.enable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(2700));
        #1us;
    endtask
endclass

class brt_usb_sof_crc5err_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_sof_crc5err_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_sof_crc5err_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        // Change ERROR to WARNING
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 1024;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 1024;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (                          ) // = 'hff
                             ,.epnum         (                          ) // = 'h1f
                             ,.dir           (                          ) // = 'b11
                             ,.pid           (  brt_usb_packet::SOF     ) // = brt_usb_packet::EXT
                             ,.crc5_err      (  1                       ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (                          ) // = 'hff
                                     ,.epnum         (                          ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::SOF     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (  1                       ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (                          ) // = 'b11
                                     );
        
        isochronous_out_xfer(.set_payload_size(1011));
        isochronous_out_xfer(.set_payload_size(1004));
        #1us;
    endtask
endclass

class brt_usb_iso_out_mps512_token_pid_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_mps512_token_pid_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_mps512_token_pid_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 512;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 512;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  4                       ) // = 'h1f
                                     ,.dir           (  0                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (  1                       ) // = 'b11
                                     ,.crc5_err      (                          ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(300));
        //mult_sb.enable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(300));
        #1us;
    endtask
endclass

class brt_usb_iso_out_mps512_token_crc5_vseq extends brt_usb_base_virtual_sequence;

    `uvm_object_utils_begin(brt_usb_iso_out_mps512_token_crc5_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_out_mps512_token_crc5_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));
        host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_FATAL),.id("DEV_CHK_TOKEN"),.new_severity(UVM_WARNING));
        //dev_agt.ulayer.link_mon.set_report_severity_override(.cur_severity(UVM_ERROR),.new_severity(UVM_WARNING));
        dev_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_override(.cur_severity(UVM_FATAL),.new_severity(UVM_WARNING));
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 512;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 512;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  4                       ) // = 'h1f
                             ,.dir           (  0                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (                          ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        host_util_cb.add_inject_err (
                                      .addr          (  0                       ) // = 'hff
                                     ,.epnum         (  4                       ) // = 'h1f
                                     ,.dir           (  0                       ) // = 'b11
                                     ,.pid           (  brt_usb_packet::OUT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     ,.pkt_err       (                          ) // = 'b00
                                     ,.pid_err       (                          ) // = 'b11
                                     ,.crc5_err      (  1                       ) // = 'b11
                                     ,.crc16_err     (                          ) // = 'b11
                                     ,.bit_stuff_err (                          ) // = 'b11
                                     ,.need_timeout  (  1                       ) // = 'b11
                                     );
        
        mult_sb.disable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(300));
        //mult_sb.enable_sb (4,0);                                         
        isochronous_out_xfer(.set_payload_size(300));
        #1us;
    endtask
endclass

// LPM protocol
class brt_usb_lpm_normal_vseq extends brt_usb_base_virtual_sequence;
    bit                                             pass;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;

    `uvm_object_utils_begin(brt_usb_lpm_normal_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_lpm_normal_vseq");
        super.new(name);
    endfunction

    virtual task body();
        super.body();
        // Change config
        host_cfg.remote_device_cfg[0].device_address = 127;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        fork
            // CTRL
            begin
                // Checker
                chk_pkt = new("chk_pkt", host_util_cb);
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA0   ) // DATA0 is same value with LPM
                                     ,.data_size     (                          ) // = -1
                                     );
                host_util_cb.add_chk_pkt(chk_pkt);

                lpm_xfer (.remote_wake(1), .hird(10), .link_state(2), .pass(pass));
                #100us;
                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;

                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                lpm_xfer (.remote_wake(1), .hird(2), .link_state(2), .pass(pass));

                #100us;

                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;
            end
        join
    endtask

    task lpm_xfer (bit remote_wake, bit [3:0] hird, bit [3:0] link_state, output bit pass);
        brt_usb_lpm_xfer_sequence  lpm_seq;
        fork
            begin
                lpm_seq = new ();
                lpm_seq.randomize() with { seq_remote_wake == remote_wake;
                                           seq_hird        == hird;
                                           seq_link_state  == link_state;
                                             };
                lpm_seq.start (p_sequencer.xfer_sequencer);
                `brt_info(get_name(), $sformatf("Done %s transfer, EP: %d", lpm_seq.req.xfer_type.name(), lpm_seq.req.endpoint_number), UVM_LOW)
                // return result
                pass = lpm_seq.req.tfer_status == brt_usb_types::ACCEPT;
            end
        join
    endtask:lpm_xfer
endclass

class brt_usb_lpm_dev_resume_vseq extends brt_usb_base_virtual_sequence;
    bit                                             pass;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;

    `uvm_object_utils_begin(brt_usb_lpm_dev_resume_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_lpm_dev_resume_vseq");
        super.new(name);
    endfunction

    virtual task body();
        super.body();
        // Change config
        host_cfg.remote_device_cfg[0].device_address = 127;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        fork
            // CTRL
            begin
                // Checker
                chk_pkt = new("chk_pkt", host_util_cb);
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA0   ) // DATA0 is same value with LPM
                                     ,.data_size     (                          ) // = -1
                                     );
                host_util_cb.add_chk_pkt(chk_pkt);

                lpm_xfer (.remote_wake(1), .hird(10), .link_state(2), .pass(pass));
                #100us;
                // Dev resume
                `brt_do_on(resume_seq, dev_agt.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;

                // Dev resume
                `brt_do_on(resume_seq, dev_agt.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                lpm_xfer (.remote_wake(1), .hird(2), .link_state(2), .pass(pass));

                #100us;

                // Dev resume
                `brt_do_on(resume_seq, dev_agt.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;
            end
        join
    endtask

    task lpm_xfer (bit remote_wake, bit [3:0] hird, bit [3:0] link_state, output bit pass);
        brt_usb_lpm_xfer_sequence  lpm_seq;
        fork
            begin
                lpm_seq = new ();
                lpm_seq.randomize() with { seq_remote_wake == remote_wake;
                                           seq_hird        == hird;
                                           seq_link_state  == link_state;
                                             };
                lpm_seq.start (p_sequencer.xfer_sequencer);
                `brt_info(get_name(), $sformatf("Done %s transfer, EP: %d", lpm_seq.req.xfer_type.name(), lpm_seq.req.endpoint_number), UVM_LOW)
                // return result
                pass = lpm_seq.req.tfer_status == brt_usb_types::ACCEPT;
            end
        join
    endtask:lpm_xfer
endclass

class brt_usb_lpm_nyet_vseq extends brt_usb_base_virtual_sequence;
    bit                                             pass;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;

    `uvm_object_utils_begin(brt_usb_lpm_nyet_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_lpm_nyet_vseq");
        super.new(name);
    endfunction

    virtual task body();
        super.body();
        // Change config
        host_cfg.remote_device_cfg[0].device_address = 127;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        fork
            // CTRL
            begin
                // Checker
                chk_pkt = new("chk_pkt", host_util_cb);
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA0   ) // DATA0 is same value with LPM
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::NYET    ) // 
                                     ,.data_size     (                          ) // = -1
                                     );
                host_util_cb.add_chk_pkt(chk_pkt);
                // error injection
                dev_util_cb.add_inject_err (
                                              .addr          (  127                     ) // = 'hff
                                             ,.epnum         (  0                       ) // = 'h1f
                                             ,.dir           (                          ) // = 'b11
                                             ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                             ,.new_pid       (  brt_usb_packet::NYET    ) // = brt_usb_packet::EXT
                                             ,.ack_pkt       (  1                       ) // = ACK of LPM transfer
                                             ,.pkt_err       (                          ) // = 'b00
                                             ,.pid_err       (                          ) // = 'b11
                                             ,.crc5_err      (                          ) // = 'b11
                                             ,.crc16_err     (                          ) // = 'b11
                                             ,.bit_stuff_err (                          ) // = 'b11
                                             ,.need_timeout  (                          ) // = 'b11
                                             ,.pkt_idx       (                          ) // = -1
                                             );

                lpm_xfer (.remote_wake(1), .hird(10), .link_state(2), .pass(pass));
                #100us;
                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #100us;
                lpm_xfer (.remote_wake(1), .hird(2), .link_state(2), .pass(pass));

                #100us;

                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;
            end
        join
    endtask

    task lpm_xfer (bit remote_wake, bit [3:0] hird, bit [3:0] link_state, output bit pass);
        brt_usb_lpm_xfer_sequence  lpm_seq;
        fork
            begin
                lpm_seq = new ();
                lpm_seq.randomize() with { seq_remote_wake == remote_wake;
                                           seq_hird        == hird;
                                           seq_link_state  == link_state;
                                             };
                lpm_seq.start (p_sequencer.xfer_sequencer);
                `brt_info(get_name(), $sformatf("Done %s transfer, EP: %d", lpm_seq.req.xfer_type.name(), lpm_seq.req.endpoint_number), UVM_LOW)
                // return result
                pass = lpm_seq.req.tfer_status == brt_usb_types::ACCEPT;
            end
        join
    endtask:lpm_xfer
endclass

class brt_usb_lpm_stall_vseq extends brt_usb_base_virtual_sequence;
    bit                                             pass;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;

    `uvm_object_utils_begin(brt_usb_lpm_stall_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_lpm_stall_vseq");
        super.new(name);
    endfunction

    virtual task body();
        super.body();
        // Change config
        host_cfg.remote_device_cfg[0].device_address = 127;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        fork
            // CTRL
            begin
                // Checker
                chk_pkt = new("chk_pkt", host_util_cb);
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA0   ) // DATA0 is same value with LPM
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::STALL   ) // 
                                     ,.data_size     (                          ) // = -1
                                     );
                host_util_cb.add_chk_pkt(chk_pkt);
                // error injection
                dev_util_cb.add_inject_err (
                                              .addr          (  127                     ) // = 'hff
                                             ,.epnum         (  0                       ) // = 'h1f
                                             ,.dir           (                          ) // = 'b11
                                             ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                             ,.new_pid       (  brt_usb_packet::STALL   ) // = brt_usb_packet::EXT
                                             ,.ack_pkt       (  1                       ) // = ACK of LPM transfer
                                             ,.pkt_err       (                          ) // = 'b00
                                             ,.pid_err       (                          ) // = 'b11
                                             ,.crc5_err      (                          ) // = 'b11
                                             ,.crc16_err     (                          ) // = 'b11
                                             ,.bit_stuff_err (                          ) // = 'b11
                                             ,.need_timeout  (                          ) // = 'b11
                                             ,.pkt_idx       (                          ) // = -1
                                             );

                lpm_xfer (.remote_wake(1), .hird(1), .link_state(2), .pass(pass));

                #1ms;
                lpm_xfer (.remote_wake(1), .hird(2), .link_state(2), .pass(pass));

                #100us;

                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;
            end
        join
    endtask

    task lpm_xfer (bit remote_wake, bit [3:0] hird, bit [3:0] link_state, output bit pass);
        brt_usb_lpm_xfer_sequence  lpm_seq;
        fork
            begin
                lpm_seq = new ();
                lpm_seq.randomize() with { seq_remote_wake == remote_wake;
                                           seq_hird        == hird;
                                           seq_link_state  == link_state;
                                             };
                lpm_seq.start (p_sequencer.xfer_sequencer);
                `brt_info(get_name(), $sformatf("Done %s transfer, EP: %d", lpm_seq.req.xfer_type.name(), lpm_seq.req.endpoint_number), UVM_LOW)
                // return result
                pass = lpm_seq.req.tfer_status == brt_usb_types::ACCEPT;
            end
        join
    endtask:lpm_xfer
endclass

class brt_usb_lpm_timeout_vseq extends brt_usb_base_virtual_sequence;
    bit                                             pass;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;

    `uvm_object_utils_begin(brt_usb_lpm_timeout_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_lpm_timeout_vseq");
        super.new(name);
    endfunction

    virtual task body();
        super.body();
        // Change config
        host_cfg.remote_device_cfg[0].device_address = 127;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        fork
            // CTRL
            begin
                // Checker
                chk_pkt = new("chk_pkt", host_util_cb);
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA0   ) // DATA0 is same value with LPM
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                host_util_cb.add_chk_pkt(chk_pkt);
                // error injection
                host_util_cb.add_inject_err (
                                              .addr          (  127                     ) // = 'hff
                                             ,.epnum         (  0                       ) // = 'h1f
                                             ,.dir           (                          ) // = 'b11
                                             ,.pid           (                          ) // = brt_usb_packet::EXT
                                             ,.lpm_pkt       (  1                       ) // = ACK of LPM transfer
                                             ,.pkt_err       (                          ) // = 'b00
                                             ,.pid_err       (                          ) // = 'b11
                                             ,.crc5_err      (                          ) // = 'b11
                                             ,.crc16_err     (                          ) // = 'b11
                                             ,.drop          (                          ) // = 'b11
                                             ,.need_timeout  (  1                       ) // = 'b11
                                             ,.pkt_idx       (                          ) // = -1
                                             );
                dev_util_cb.add_inject_err (
                                              .addr          (  127                     ) // = 'hff
                                             ,.epnum         (  0                       ) // = 'h1f
                                             ,.dir           (                          ) // = 'b11
                                             ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                             ,.ack_pkt       (  1                       ) // = ACK of LPM transfer
                                             ,.pkt_err       (                          ) // = 'b00
                                             ,.pid_err       (                          ) // = 'b11
                                             ,.crc5_err      (                          ) // = 'b11
                                             ,.crc16_err     (                          ) // = 'b11
                                             ,.drop          (  1                         ) // = 'b11
                                             ,.need_timeout  (                          ) // = 'b11
                                             ,.pkt_idx       (                          ) // = -1
                                             );

                lpm_xfer (.remote_wake(1), .hird(1), .link_state(2), .pass(pass));

                #100us;
                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #1ms;
                lpm_xfer (.remote_wake(1), .hird(2), .link_state(2), .pass(pass));

                #100us;

                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;
            end
        join
    endtask

    task lpm_xfer (bit remote_wake, bit [3:0] hird, bit [3:0] link_state, output bit pass);
        brt_usb_lpm_xfer_sequence  lpm_seq;
        fork
            begin
                lpm_seq = new ();
                lpm_seq.randomize() with { seq_remote_wake == remote_wake;
                                           seq_hird        == hird;
                                           seq_link_state  == link_state;
                                             };
                lpm_seq.start (p_sequencer.xfer_sequencer);
                `brt_info(get_name(), $sformatf("Done %s transfer, EP: %d", lpm_seq.req.xfer_type.name(), lpm_seq.req.endpoint_number), UVM_LOW)
                // return result
                pass = lpm_seq.req.tfer_status == brt_usb_types::ACCEPT;
            end
        join
    endtask:lpm_xfer
endclass

class brt_usb_lpm_ack_piderr_vseq extends brt_usb_base_virtual_sequence;
    bit                                             pass;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;

    `uvm_object_utils_begin(brt_usb_lpm_ack_piderr_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_lpm_ack_piderr_vseq");
        super.new(name);
    endfunction

    virtual task body();
        super.body();
        // Change config
        host_cfg.remote_device_cfg[0].device_address = 127;
        // disable monitor checker
        host_cfg.ignore_mon_host_err = 1;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        fork
            // CTRL
            begin
                // Checker
                chk_pkt = new("chk_pkt", host_util_cb);
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::DATA0   ) // DATA0 is same value with LPM
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                host_util_cb.add_chk_pkt(chk_pkt);
                // error injection
                host_util_cb.add_inject_err (
                                              .addr          (  127                     ) // = 'hff
                                             ,.epnum         (  0                       ) // = 'h1f
                                             ,.dir           (                          ) // = 'b11
                                             ,.pid           (                          ) // = brt_usb_packet::EXT
                                             ,.lpm_pkt       (  1                       ) // = ACK of LPM transfer
                                             ,.pkt_err       (                          ) // = 'b00
                                             ,.pid_err       (                          ) // = 'b11
                                             ,.crc5_err      (                          ) // = 'b11
                                             ,.crc16_err     (                          ) // = 'b11
                                             ,.drop          (                          ) // = 'b11
                                             ,.need_timeout  (                          ) // = 'b11
                                             ,.pkt_idx       (                          ) // = -1
                                             );
                dev_util_cb.add_inject_err (
                                              .addr          (  127                     ) // = 'hff
                                             ,.epnum         (  0                       ) // = 'h1f
                                             ,.dir           (                          ) // = 'b11
                                             ,.pid           (  brt_usb_packet::ACK     ) // = brt_usb_packet::EXT
                                             ,.ack_pkt       (  1                       ) // = ACK of LPM transfer
                                             ,.pkt_err       (                          ) // = 'b00
                                             ,.pid_err       (  1                       ) // = 'b11
                                             ,.crc5_err      (                          ) // = 'b11
                                             ,.crc16_err     (                          ) // = 'b11
                                             ,.drop          (                            ) // = 'b11
                                             ,.need_timeout  (                          ) // = 'b11
                                             ,.pkt_idx       (                          ) // = -1
                                             );

                lpm_xfer (.remote_wake(1), .hird(1), .link_state(2), .pass(pass));

                #100us;
                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #1ms;
                lpm_xfer (.remote_wake(1), .hird(2), .link_state(2), .pass(pass));

                #100us;

                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;
            end
        join
    endtask

    task lpm_xfer (bit remote_wake, bit [3:0] hird, bit [3:0] link_state, output bit pass);
        brt_usb_lpm_xfer_sequence  lpm_seq;
        fork
            begin
                lpm_seq = new ();
                lpm_seq.randomize() with { seq_remote_wake == remote_wake;
                                           seq_hird        == hird;
                                           seq_link_state  == link_state;
                                             };
                lpm_seq.start (p_sequencer.xfer_sequencer);
                `brt_info(get_name(), $sformatf("Done %s transfer, EP: %d", lpm_seq.req.xfer_type.name(), lpm_seq.req.endpoint_number), UVM_LOW)
                // return result
                pass = lpm_seq.req.tfer_status == brt_usb_types::ACCEPT;
            end
        join
    endtask:lpm_xfer
endclass

class brt_usb_lpm_ack_exterr_lpmerr_vseq extends brt_usb_base_virtual_sequence;
    bit                                             pass;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;

    `uvm_object_utils_begin(brt_usb_lpm_ack_exterr_lpmerr_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_lpm_ack_exterr_lpmerr_vseq");
        super.new(name);
    endfunction

    virtual task body();
        super.body();
        // Change config
        host_cfg.remote_device_cfg[0].device_address = 127;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        fork
            // CTRL
            begin
                // Checker
                chk_pkt = new("chk_pkt", host_util_cb);
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.pid_err       (  1                       ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                chk_pkt.add_chk_pnt (
                                      .addr          (  127                     ) // = 'hff
                                     ,.epnum         (  0                       ) // = 'h1f
                                     ,.dir           (                          ) // = 'b11
                                     ,.pid           (  brt_usb_packet::EXT     ) // = brt_usb_packet::EXT
                                     ,.data_size     (                          ) // = -1
                                     );
                host_util_cb.add_chk_pkt(chk_pkt);
                // error injection
                host_util_cb.add_inject_err (
                                              .addr          (  127                     ) // = 'hff
                                             ,.epnum         (  0                       ) // = 'h1f
                                             ,.dir           (                          ) // = 'b11
                                             ,.pid           (                          ) // = brt_usb_packet::EXT
                                             ,.ext_pkt       (  1                       ) // = ACK of LPM transfer
                                             ,.pkt_err       (                          ) // = 'b00
                                             ,.pid_err       (  1                       ) // = 'b11
                                             ,.crc5_err      (                          ) // = 'b11
                                             ,.crc16_err     (                          ) // = 'b11
                                             ,.drop          (                          ) // = 'b11
                                             ,.need_timeout  (                          ) // = 'b11
                                             ,.pkt_idx       (                          ) // = -1
                                             );
                host_util_cb.add_inject_err (
                                              .addr          (  127                     ) // = 'hff
                                             ,.epnum         (  0                       ) // = 'h1f
                                             ,.dir           (                          ) // = 'b11
                                             ,.pid           (                          ) // = brt_usb_packet::EXT
                                             ,.lpm_pkt       (  1                       ) // = ACK of LPM transfer
                                             ,.pkt_err       (                          ) // = 'b00
                                             ,.pid_err       (  1                       ) // = 'b11
                                             ,.crc5_err      (                          ) // = 'b11
                                             ,.crc16_err     (                          ) // = 'b11
                                             ,.drop          (                          ) // = 'b11
                                             ,.need_timeout  (  1                       ) // = 'b11
                                             ,.pkt_idx       (                          ) // = -1
                                             );

                lpm_xfer (.remote_wake(1), .hird(1), .link_state(2), .pass(pass));

                #100us;
                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #1ms;
                lpm_xfer (.remote_wake(1), .hird(2), .link_state(2), .pass(pass));

                #100us;

                // Host resume
                `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
                wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

                #10ms;
            end
        join
    endtask

    task lpm_xfer (bit remote_wake, bit [3:0] hird, bit [3:0] link_state, output bit pass);
        brt_usb_lpm_xfer_sequence  lpm_seq;
        fork
            begin
                lpm_seq = new ();
                lpm_seq.randomize() with { seq_remote_wake == remote_wake;
                                           seq_hird        == hird;
                                           seq_link_state  == link_state;
                                             };
                lpm_seq.start (p_sequencer.xfer_sequencer);
                `brt_info(get_name(), $sformatf("Done %s transfer, EP: %d", lpm_seq.req.xfer_type.name(), lpm_seq.req.endpoint_number), UVM_LOW)
                // return result
                pass = lpm_seq.req.tfer_status == brt_usb_types::ACCEPT;
            end
        join
    endtask:lpm_xfer
endclass

class brt_usb_iso_in_lpm_vseq extends brt_usb_base_virtual_sequence;
    bit                                             pass;
    brt_usb_link_service_clear_suspend_sequence     resume_seq;

    `uvm_object_utils_begin(brt_usb_iso_in_lpm_vseq)
    `uvm_object_utils_end

    function new(string name="brt_usb_iso_in_lpm_vseq");
        super.new(name);
        //err_inject_cb = new();
    endfunction

    virtual task body();
        super.body();
        init_callback();
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[3].max_packet_size = 77;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_burst_size  = 0;
        p_sequencer.agt.cfg.remote_device_cfg[0].endpoint_cfg[4].max_packet_size = 77;
        reset_dev();
        start_xfer();
    endtask

    virtual task start_xfer();
        brt_usb_protocol_service_20_sof_on_off_sequence     sof_seq;

        brt_usb_base_control_xfer_sequence ctrl_seq;

        // Change ERROR to WARNING
        //host_agt.ulayer.brt_usb_20_pkt_sequencer.set_report_severity_id_override(.cur_severity(UVM_ERROR),.id("EP_BW"),.new_severity(UVM_WARNING));

        // Start SOF
        `uvm_info(get_name(), $sformatf("Start SOF"), UVM_LOW)
        `uvm_do_on_with(sof_seq, p_sequencer.prot_service_sequencer, {sof_on == 1;}) 
        `uvm_info(get_name(), $sformatf("Done starting SOF"), UVM_LOW)

        // Checker
        chk_pkt = new("chk_pkt", host_util_cb);
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  77                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        chk_pkt.add_chk_pnt (
                              .addr          (  0                       ) // = 'hff
                             ,.epnum         (  3                       ) // = 'h1f
                             ,.dir           (  1                       ) // = 'b11
                             ,.pid           (  brt_usb_packet::DATA0   ) // = brt_usb_packet::EXT
                             ,.data_size     (  55                      ) // = -1
                             ,.pkt_idx       (                          ) // = -1
                             );
        host_util_cb.add_chk_pkt(chk_pkt);
        
        isochronous_in_xfer(.set_payload_size(77));
        lpm_xfer (.remote_wake(1), .hird(1), .link_state(2), .pass(pass));

        #700us;
        // Host resume
        `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
        wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

        isochronous_in_xfer(.set_payload_size(55));
        lpm_xfer (.remote_wake(1), .hird(1), .link_state(2), .pass(pass));

        #700us;
        // Host resume
        `brt_do_on(resume_seq, p_sequencer.link_service_sequencer) 
        wait (p_sequencer.link_service_sequencer.agt.shared_status.link_usb_20_state == brt_usb_types::ENABLED);

        isochronous_in_xfer(.set_payload_size(44));
    endtask

    task lpm_xfer (bit remote_wake, bit [3:0] hird, bit [3:0] link_state, output bit pass);
        brt_usb_lpm_xfer_sequence  lpm_seq;
        fork
            begin
                lpm_seq = new ();
                lpm_seq.randomize() with { seq_remote_wake == remote_wake;
                                           seq_hird        == hird;
                                           seq_link_state  == link_state;
                                             };
                lpm_seq.start (p_sequencer.xfer_sequencer);
                `brt_info(get_name(), $sformatf("Done %s transfer, EP: %d", lpm_seq.req.xfer_type.name(), lpm_seq.req.endpoint_number), UVM_LOW)
                // return result
                pass = lpm_seq.req.tfer_status == brt_usb_types::ACCEPT;
            end
        join
    endtask:lpm_xfer
endclass