package brt_usb_env_pkg;

`include "brt_uvm_methodology.svh"

import brt_usb_pkg::*;

`include "brt_usb_scoreboard.sv"
`include "brt_usb_env.sv"

endpackage
