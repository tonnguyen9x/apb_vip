package brt_usb_pkg;
  `include "brt_usb_timescale.sv"

typedef class brt_usb_agent;

  `include "brt_uvm_methodology.svh"
  `include "brt_usb_defs.svh"
  `include "brt_usb_types.sv"
  `include "brt_usb_base_config.sv"
  `include "brt_usb_transfer.sv"
  `include "brt_usb_service.sv"
  `include "brt_usb_sequencer.sv"
  `include "brt_usb_monitor.sv"
  `include "brt_usb_base_seq_lib.sv"
  `include "brt_usb_dev_reactive.sv"
  `include "brt_usb_layering.sv"
  `include "brt_usb_driver.sv"
  `include "brt_usb_cov_wrapper.sv"
  `include "brt_usb_callbacks.sv"
  `include "brt_usb_agent.sv"

endpackage
