timeunit 1ps;
timeprecision 1ps;
