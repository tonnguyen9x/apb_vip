`include "brt_usb_protocol_service_20_sof_on_off_sequence.svh"
`include "brt_usb_packet_base_sequence.svh"
`include "brt_usb_virtual_sequence.svh"
`include "brt_usb_packet2data_sequence.svh"
`include "brt_usb_xfer2packet_sequence.svh"
`include "brt_usb_sof_pkt_sequence.svh"
`include "brt_usb_protservice_sequence.svh"
`include "brt_usb_linkservice_sequence.svh"
`include "brt_usb_link_service_packet_sequence.svh"
`include "brt_usb_device_response_sequence.svh"
`include "brt_usb_agent_wait_for_link_usb_20_state_virtual_sequence.svh"
`include "brt_usb_xfer_router_sequence.svh"
`include "brt_usb_xfer_base_sequence.svh"
`include "brt_usb_lpm_xfer_sequence.svh"
`include "brt_usb_bad_packet.svh"
