`include "brt_usb_base_control_xfer_sequence.sv"

`include "brt_usb_base_random_xfer_sequence.sv"
`include "brt_usb_base_bulk_in_xfer_sequence.sv"
`include "brt_usb_base_bulk_out_xfer_sequence.sv"

`include "brt_usb_base_interrupt_in_xfer_sequence.sv"
`include "brt_usb_base_interrupt_out_xfer_sequence.sv"

`include "brt_usb_base_random_isochronous_xfer_sequence.sv"
`include "brt_usb_base_isochronous_in_xfer_sequence.sv"
`include "brt_usb_base_isochronous_out_xfer_sequence.sv"

//`include "enumeration_sequence.sv"
//`include "enum_bulk_out_sequence.sv"
//`include "enum_bulk_in_sequence.sv"
//`include "enum_interrupt_out_sequence.sv"
//`include "enum_interrupt_in_sequence.sv"
//`include "enum_isochronous_out_sequence.sv"
//`include "enum_isochronous_in_sequence.sv"
//`include "enum_bulk_loopback.sv"
//
//`include "nyet_ping_sequence.sv"
//`include "random_data_ready_sequence.sv"
//`include "random_nak_sequence.sv"
//`include "random_stall_sequence.sv"
//`include "bad_address_sequence.sv"
//
//`include "reset_handshake_sequence.sv"
